module adc (clk,
    ready,
    start,
    analog_in,
    data_out);
 input clk;
 output ready;
 input start;
 input [7:0] analog_in;
 output [7:0] data_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net9;
 wire net19;
 wire net;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;

 sg13g2_mux2_1 _17_ (.A0(net35),
    .A1(net1),
    .S(net19),
    .X(_05_));
 sg13g2_mux2_1 _18_ (.A0(net33),
    .A1(net2),
    .S(net19),
    .X(_06_));
 sg13g2_mux2_1 _19_ (.A0(net29),
    .A1(net3),
    .S(net19),
    .X(_07_));
 sg13g2_mux2_1 _20_ (.A0(net34),
    .A1(net4),
    .S(net19),
    .X(_00_));
 sg13g2_mux2_1 _21_ (.A0(net32),
    .A1(net5),
    .S(net19),
    .X(_01_));
 sg13g2_mux2_1 _22_ (.A0(net30),
    .A1(net6),
    .S(net19),
    .X(_02_));
 sg13g2_mux2_1 _23_ (.A0(net31),
    .A1(net7),
    .S(net19),
    .X(_03_));
 sg13g2_mux2_1 _24_ (.A0(net28),
    .A1(net8),
    .S(net19),
    .X(_04_));
 sg13g2_dfrbpq_1 _25_ (.RESET_B(net27),
    .D(_05_),
    .Q(net10),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _26_ (.RESET_B(net26),
    .D(_06_),
    .Q(net11),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _27_ (.RESET_B(net25),
    .D(_07_),
    .Q(net12),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _28_ (.RESET_B(net24),
    .D(_00_),
    .Q(net13),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _29_ (.RESET_B(net23),
    .D(_01_),
    .Q(net14),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _30_ (.RESET_B(net22),
    .D(_02_),
    .Q(net15),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _31_ (.RESET_B(net21),
    .D(_03_),
    .Q(net16),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _32_ (.RESET_B(net),
    .D(_04_),
    .Q(net17),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _33_ (.RESET_B(net20),
    .D(net9),
    .Q(net18),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_tiehi _33__21 (.L_HI(net20));
 sg13g2_tiehi _31__22 (.L_HI(net21));
 sg13g2_tiehi _30__23 (.L_HI(net22));
 sg13g2_tiehi _29__24 (.L_HI(net23));
 sg13g2_tiehi _28__25 (.L_HI(net24));
 sg13g2_tiehi _27__26 (.L_HI(net25));
 sg13g2_tiehi _26__27 (.L_HI(net26));
 sg13g2_tiehi _25__28 (.L_HI(net27));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_1 input1 (.A(analog_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(analog_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(analog_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(analog_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(analog_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(analog_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(analog_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(analog_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(start),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(data_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(data_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(data_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(data_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(data_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(data_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(data_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(data_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(ready));
 sg13g2_buf_1 fanout19 (.A(net9),
    .X(net19));
 sg13g2_tiehi _32__20 (.L_HI(net));
 sg13g2_buf_16 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold29 (.A(net17),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold30 (.A(net12),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold31 (.A(net15),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold32 (.A(net16),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold33 (.A(net14),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold34 (.A(net11),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold35 (.A(net13),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold36 (.A(net10),
    .X(net35));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_fill_2 FILLER_0_42 ();
 sg13g2_fill_1 FILLER_0_44 ();
 sg13g2_decap_8 FILLER_0_53 ();
 sg13g2_fill_2 FILLER_0_60 ();
 sg13g2_fill_1 FILLER_0_62 ();
 sg13g2_decap_8 FILLER_0_71 ();
 sg13g2_decap_8 FILLER_0_78 ();
 sg13g2_decap_8 FILLER_0_85 ();
 sg13g2_decap_8 FILLER_0_92 ();
 sg13g2_fill_2 FILLER_0_99 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_67 ();
 sg13g2_decap_8 FILLER_1_74 ();
 sg13g2_decap_8 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_102 ();
 sg13g2_decap_8 FILLER_1_109 ();
 sg13g2_decap_8 FILLER_1_116 ();
 sg13g2_decap_8 FILLER_1_123 ();
 sg13g2_decap_8 FILLER_1_130 ();
 sg13g2_decap_8 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_fill_1 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_1 FILLER_3_52 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_4 FILLER_4_42 ();
 sg13g2_fill_2 FILLER_4_46 ();
 sg13g2_decap_4 FILLER_4_52 ();
 sg13g2_fill_2 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_72 ();
 sg13g2_decap_8 FILLER_4_82 ();
 sg13g2_decap_8 FILLER_4_89 ();
 sg13g2_decap_4 FILLER_4_96 ();
 sg13g2_fill_2 FILLER_4_100 ();
 sg13g2_fill_2 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_118 ();
 sg13g2_fill_1 FILLER_4_120 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_fill_2 FILLER_4_151 ();
 sg13g2_fill_1 FILLER_4_153 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_4 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_136 ();
 sg13g2_decap_8 FILLER_5_143 ();
 sg13g2_decap_4 FILLER_5_150 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_decap_4 FILLER_6_141 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_127 ();
 sg13g2_decap_8 FILLER_7_134 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_decap_4 FILLER_7_148 ();
 sg13g2_fill_2 FILLER_7_152 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_131 ();
 sg13g2_decap_8 FILLER_8_142 ();
 sg13g2_decap_4 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_fill_2 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_31 ();
 sg13g2_fill_1 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_45 ();
 sg13g2_decap_8 FILLER_10_52 ();
 sg13g2_decap_8 FILLER_10_59 ();
 sg13g2_decap_8 FILLER_10_66 ();
 sg13g2_decap_8 FILLER_10_73 ();
 sg13g2_decap_8 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_87 ();
 sg13g2_decap_8 FILLER_10_94 ();
 sg13g2_decap_8 FILLER_10_101 ();
 sg13g2_decap_8 FILLER_10_108 ();
 sg13g2_decap_4 FILLER_10_115 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_4 FILLER_10_144 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_decap_8 FILLER_11_8 ();
 sg13g2_decap_4 FILLER_11_15 ();
 sg13g2_fill_1 FILLER_11_19 ();
 sg13g2_decap_8 FILLER_11_47 ();
 sg13g2_decap_8 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_decap_8 FILLER_11_75 ();
 sg13g2_decap_8 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_89 ();
 sg13g2_decap_8 FILLER_11_96 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_8 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_29 ();
 sg13g2_decap_8 FILLER_12_36 ();
 sg13g2_decap_8 FILLER_12_43 ();
 sg13g2_decap_8 FILLER_12_50 ();
 sg13g2_decap_8 FILLER_12_57 ();
 sg13g2_decap_8 FILLER_12_64 ();
 sg13g2_decap_8 FILLER_12_71 ();
 sg13g2_decap_8 FILLER_12_78 ();
 sg13g2_decap_8 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_decap_8 FILLER_12_99 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_117 ();
 sg13g2_decap_8 FILLER_12_124 ();
 sg13g2_decap_8 FILLER_12_131 ();
 sg13g2_decap_8 FILLER_12_138 ();
 sg13g2_decap_8 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_fill_2 FILLER_13_25 ();
 sg13g2_fill_1 FILLER_13_27 ();
 sg13g2_decap_4 FILLER_13_38 ();
 sg13g2_fill_2 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_decap_8 FILLER_13_71 ();
 sg13g2_decap_8 FILLER_13_78 ();
 sg13g2_decap_8 FILLER_13_85 ();
 sg13g2_decap_4 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_decap_8 FILLER_13_135 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_4 FILLER_14_25 ();
 sg13g2_decap_4 FILLER_14_33 ();
 sg13g2_decap_8 FILLER_14_64 ();
 sg13g2_decap_4 FILLER_14_71 ();
 sg13g2_decap_4 FILLER_14_113 ();
 sg13g2_fill_1 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_127 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_decap_4 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_decap_4 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_152 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_4 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_100 ();
 sg13g2_decap_8 FILLER_16_107 ();
 sg13g2_decap_8 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_121 ();
 sg13g2_decap_8 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_135 ();
 sg13g2_decap_8 FILLER_16_142 ();
 sg13g2_decap_4 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_69 ();
 sg13g2_decap_8 FILLER_18_76 ();
 sg13g2_decap_8 FILLER_18_83 ();
 sg13g2_decap_8 FILLER_18_90 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_117 ();
 sg13g2_decap_8 FILLER_18_124 ();
 sg13g2_decap_8 FILLER_18_131 ();
 sg13g2_decap_8 FILLER_18_138 ();
 sg13g2_decap_8 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_152 ();
endmodule
